/******************************************************************************
Author: Hyoukjun Kwon (hyoukjun@gatech.edu)

Copyright (c) 2017 Georgia Instititue of Technology

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
SOFTWARE.

*******************************************************************************/

/* Primitives */
import Vector::*;

/* Microswitch types */
import MicroswitchTypes::*;
import MicroswitchMessageTypes::*;

/* Neural network types */
import NeuralNetworkConfig::*;
import NeuralNetworkTypes::*;

//Assumption: NumPEs = 2^n
typedef TLog#(NumPEs)                          MS_NumMicroswitchLevels;
typedef MS_NumMicroswitchLevels                MS_NumMiddleSwitchLevels;
typedef TMul#(MS_NumMicroswitchLevels, NumPEs) MS_NumSwitches; // N log(N)
typedef TDiv#(NumPEs, 2)                       MS_NumLowestBranchNodes;
typedef TSub#(NumPEs, 1)                       MS_NumBranchNodes; // N-1

typedef TDiv#(NumPEs, 2)                       MS_RootTopSwitchID;

interface NetworkExternalInterface;
  method Action putFlit(Flit req);
  method ActionValue#(Flit) getFlit;
endinterface

typedef Vector#(MS_NumBranchNodes, MS_SetupSignal) MS_ScatterSetupSignal;
